module d_ff_tb();
 reg d0, d1,sel,rstclk;
 wire q;
 
 // Module Instantiation
 dff DUT()
 
    
  
