module d_ff_tb();
 
    
  
